module RAM;

logic[7:0] core[256];

endmodule