module ROM;

logic[8:0] core[65536];

endmodule